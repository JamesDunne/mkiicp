****************************************************
.SUBCKT 12AX7 1 2 3; A G C;
*      Extract V3.000
* Model created: 16-Dec-2020  by kurtblum.com
*
X1 1 2 3 TriodeK MU= 96.20 EX=1.437 KG1= 613.4 KP= 740.3 KVB= 1672. RGI=2000
+ CCG=0.0P  CGP=0.0P CCP=0.0P  ;
.ENDS
 
****************************************************
.SUBCKT TriodeK 1 2 3; A G C
*
* NOTE: LOG(x) is base e LOG or natural logarithm.
* For some Spice versions, e.g. MicroCap, this has to be changed to LN(x).
*
E1 7 0 VALUE=
+{V(1,3)/KP*LOG(1+EXP(KP*(1/MU+V(2,3)/SQRT(KVB+V(1,3)*V(1,3)))))}
RE1 7 0 1G
G1 1 3 VALUE={0.5*(PWR(V(7),EX)+PWRS(V(7),EX))/KG1}
RCP 1 3 1G    ; TO AVOID FLOATING NODES IN MU-FOLLOWER
C1 2 3 {CCG}  ; CATHODE-GRID
C2 2 1 {CGP}  ; GRID-PLATE
C3 1 3 {CCP}  ; CATHODE-PLATE
D3 5 3 DX     ; FOR GRID CURRENT
R1 2 5 {RGI}  ; FOR GRID CURRENT
.MODEL DX D(IS=1N RS=1 CJO=10PF TT=1N)
.ENDS TriodeK
